magic
tech sky130A
magscale 1 2
timestamp 1752845668
<< metal3 >>
rect 1200 440 1972 608
<< metal4 >>
rect 79 647 1601 1369
rect 1279 79 1601 401
rect 1872 12 1968 1436
use sky130_fd_pr__cap_mim_m3_1_4CW8F2  sky130_fd_pr__cap_mim_m3_1_4CW8F2_0
timestamp 1752698335
transform 1 0 986 0 1 1008
box -986 -440 986 440
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1752698335
transform 1 0 1586 0 1 240
box -386 -240 386 240
<< labels >>
flabel metal4 s 1279 79 1601 401 0 FreeSans 320 0 0 0 liltop
port 2 nsew
flabel metal4 s 79 647 1601 1369 0 FreeSans 320 0 0 0 bigtop
port 1 nsew
flabel metal4 s 1872 12 1968 1436 0 FreeSans 320 90 0 0 bottom
port 0 nsew
<< end >>

magic
tech sky130A
timestamp 1752846221
<< nwell >>
rect 30 672 508 760
rect 30 476 600 672
rect 30 334 750 476
rect 30 30 1024 334
<< pdiff >>
rect 90 613 448 702
rect 90 416 540 613
rect 90 274 690 416
rect 90 91 957 274
rect 90 90 209 91
<< psubdiff >>
rect 0 773 538 790
rect 0 17 17 773
rect 521 702 538 773
rect 521 685 630 702
rect 613 506 630 685
rect 613 489 780 506
rect 763 364 780 489
rect 763 347 1054 364
rect 1037 17 1054 347
rect 0 0 1054 17
<< nsubdiff >>
rect 48 727 490 742
rect 48 63 63 727
rect 475 654 490 727
rect 475 639 582 654
rect 567 458 582 639
rect 567 443 732 458
rect 717 316 732 443
rect 717 301 1006 316
rect 991 63 1006 301
rect 48 48 1006 63
<< end >>

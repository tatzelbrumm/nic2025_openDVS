magic
tech sky130A
timestamp 1752354234
<< isosubstrate >>
rect 0 0 1200 1200
<< end >>

* SPICE3 file created from photodiode.ext - technology: sky130A

C0 cathode guard 9.60337f

magic
tech sky130A
magscale 1 2
timestamp 1752698462
<< metal4 >>
rect -1507 407 15 1129
rect -307 -161 15 161
rect 286 -228 382 1196
use sky130_fd_pr__cap_mim_m3_1_4CW8F2  sky130_fd_pr__cap_mim_m3_1_4CW8F2_0
timestamp 1752698335
transform 1 0 -600 0 1 768
box -986 -440 986 440
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1752698335
transform 1 0 0 0 1 0
box -386 -240 386 240
<< labels >>
flabel metal4 s 286 -228 382 1196 0 FreeSans 320 90 0 0 bottom
port 0 nsew
flabel metal4 s -1507 407 15 1129 0 FreeSans 320 0 0 0 bigtop
port 1 nsew
flabel metal4 s -307 -161 15 161 0 FreeSans 320 0 0 0 liltop
port 2 nsew
<< properties >>
string FIXED_BBOX -386 -240 94 240
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

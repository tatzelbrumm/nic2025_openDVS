magic
tech sky130A
magscale 1 2
timestamp 1752834577
<< error_s >>
rect 2139 1903 2227 1914
rect 2150 1891 2216 1903
rect 1981 1880 2109 1881
rect 2139 1880 2227 1891
rect 1836 1368 1870 1415
rect 1708 1318 1779 1320
rect 1862 1318 1870 1368
rect 1708 1297 1752 1318
rect 1768 1309 1779 1318
rect 1859 1307 1870 1318
rect 1708 1286 1763 1297
rect 2020 764 2139 774
rect 2020 753 2031 764
rect 2128 763 2139 764
<< poly >>
rect 2150 1918 2216 1934
rect 2150 1884 2166 1918
rect 2202 1884 2216 1918
rect 2150 1868 2216 1884
rect 2186 1748 2216 1868
rect 1702 1368 1768 1384
rect 1702 1334 1718 1368
rect 1752 1334 1768 1368
rect 1702 1318 1768 1334
rect 1862 1368 1928 1384
rect 1862 1334 1878 1368
rect 1912 1334 1928 1368
rect 1862 1318 1928 1334
rect 1722 1230 1752 1318
rect 1898 1230 1928 1318
rect 1888 814 1954 830
rect 1888 780 1904 814
rect 1938 798 1954 814
rect 2098 798 2128 830
rect 1938 780 2128 798
rect 1888 764 2128 780
<< polycont >>
rect 2166 1884 2202 1918
rect 1718 1334 1752 1368
rect 1878 1334 1912 1368
rect 1904 780 1938 814
<< locali >>
rect 2166 2394 2202 2400
rect 1718 1962 1752 1968
rect 1718 1368 1752 1922
rect 2166 1918 2202 2354
rect 1856 1878 1892 1884
rect 2166 1868 2202 1884
rect 1856 1368 1892 1838
rect 2228 1734 2390 1752
rect 2228 1562 2354 1734
rect 2228 1544 2390 1562
rect 1856 1334 1878 1368
rect 1912 1334 1928 1368
rect 1718 1318 1752 1334
rect 1888 814 1954 830
rect 1888 780 1904 814
rect 1938 780 1954 814
rect 1888 764 1954 780
<< viali >>
rect 2166 2354 2202 2394
rect 1718 1922 1752 1962
rect 1856 1838 1892 1878
rect 2354 1562 2390 1734
rect 1904 780 1938 814
<< metal1 >>
rect 1934 1736 2100 1748
rect 1934 1560 2048 1736
rect 1934 1548 2100 1560
rect 2348 1734 2400 1746
rect 2348 1550 2400 1562
rect 2132 1482 2268 1494
rect 1030 1420 1892 1466
rect 1030 1416 1108 1420
rect 1030 1362 1042 1416
rect 1096 1362 1108 1416
rect 1030 1350 1108 1362
rect 1748 1370 1814 1388
rect 1748 1318 1754 1370
rect 1808 1318 1814 1370
rect 1748 1298 1814 1318
rect 1758 1130 1804 1298
rect 1846 1130 1892 1420
rect 2184 1306 2268 1482
rect 2132 1294 2268 1306
rect 2046 1218 2316 1230
rect 2046 842 2216 1218
rect 2046 830 2316 842
rect 1888 824 1954 830
rect 1888 770 1894 824
rect 1948 770 1954 824
rect 1888 764 1954 770
<< via1 >>
rect 1522 2132 1584 2184
rect 1754 2006 1808 2094
rect 2048 1560 2100 1736
rect 2348 1562 2354 1734
rect 2354 1562 2390 1734
rect 2390 1562 2400 1734
rect 1042 1362 1096 1416
rect 1754 1318 1808 1370
rect 2132 1306 2184 1482
rect 2216 842 2316 1218
rect 1894 814 1948 824
rect 1894 780 1904 814
rect 1904 780 1938 814
rect 1938 780 1948 814
rect 1894 770 1948 780
<< metal2 >>
rect 1518 2184 1588 2190
rect 1518 2132 1522 2184
rect 1584 2132 1588 2184
rect 1030 1418 1108 1428
rect 1030 1360 1040 1418
rect 1098 1360 1108 1418
rect 1030 1350 1108 1360
rect 1518 836 1588 2132
rect 1748 2094 1814 2100
rect 1748 2006 1754 2094
rect 1808 2006 1814 2094
rect 1748 1370 1814 2006
rect 1748 1318 1754 1370
rect 1808 1318 1814 1370
rect 1748 1312 1814 1318
rect 1514 826 1592 836
rect 1514 768 1524 826
rect 1582 768 1592 826
rect 1514 758 1592 768
rect 1872 826 1968 848
rect 1872 768 1892 826
rect 1950 768 1968 826
rect 1872 752 1968 768
<< via2 >>
rect 1040 1416 1098 1418
rect 1040 1362 1042 1416
rect 1042 1362 1096 1416
rect 1096 1362 1098 1416
rect 1040 1360 1098 1362
rect 1524 768 1582 826
rect 1892 824 1950 826
rect 1892 770 1894 824
rect 1894 770 1948 824
rect 1948 770 1950 824
rect 1892 768 1950 770
<< metal3 >>
rect 1016 1424 1120 1440
rect 1016 1356 1034 1424
rect 1104 1356 1120 1424
rect 1016 1344 1120 1356
rect 1500 832 1604 848
rect 1500 764 1518 832
rect 1588 764 1604 832
rect 1500 752 1604 764
rect 1868 832 1972 848
rect 1868 764 1886 832
rect 1956 764 1972 832
rect 1868 752 1972 764
<< via3 >>
rect 1034 1418 1104 1424
rect 1034 1360 1040 1418
rect 1040 1360 1098 1418
rect 1098 1360 1104 1418
rect 1034 1356 1104 1360
rect 1518 826 1588 832
rect 1518 768 1524 826
rect 1524 768 1582 826
rect 1582 768 1588 826
rect 1518 764 1588 768
rect 1886 826 1956 832
rect 1886 768 1892 826
rect 1892 768 1950 826
rect 1950 768 1956 826
rect 1886 764 1956 768
<< metal4 >>
rect 1020 1424 1116 1666
rect 1020 1356 1034 1424
rect 1104 1356 1116 1424
rect 1020 1344 1116 1356
rect 1504 832 1600 1072
rect 1504 764 1518 832
rect 1588 764 1600 832
rect 1504 752 1600 764
rect 1872 832 1968 964
rect 1872 764 1886 832
rect 1956 764 1968 832
rect 1872 752 1968 764
use mimcaps  mimcaps_0
timestamp 1752833958
transform 1 0 0 0 1 952
box 0 0 1972 1448
use pixeltransistors  pixeltransistors_0
timestamp 1752834206
transform 1 0 1520 0 1 1160
box 144 -420 842 754
use wires  wires_0
timestamp 1752781518
transform 1 0 0 0 1 0
box 0 0 2400 2400
<< end >>

magic
tech sky130A
timestamp 1752533151
<< metal1 >>
rect 0 14 1200 28
rect 0 42 1200 56
rect 0 70 1200 84
rect 0 1116 1200 1130
rect 0 1144 1200 1158
rect 0 1172 1200 1186
<< metal2 >>
rect 1116 0 1130 1200
rect 1144 0 1158 1200
rect 1172 0 1186 1200
<< labels >>
flabel metal1 0 14 1200 28 0 FreeSans 100 0 0 0 GND
port 0 ew
flabel metal1 0 1116 1200 1130 0 FreeSans 100 0 0 0 VDD
port 1 ew
flabel metal1 0 42 1200 56 0 FreeSans 100 0 0 0 vph_bias
port 2 ew
flabel metal1 0 70 1200 84 0 FreeSans 100 0 0 0 sf_bias
port 3 ew
flabel metal1 0 1144 1200 1158 0 FreeSans 100 0 0 0 vref
port 4 ew
flabel metal1 0 1172 1200 1186 0 FreeSans 100 0 0 0 row_sel
port 5 ew
flabel metal2 1116 0 1130 1200 0 FreeSans 100 90 0 0 sense
port 6 ns
flabel metal2 1144 0 1158 1200 0 FreeSans 100 90 0 0 feedback
port 7 ns
flabel metal2 1172 0 1186 1200 0 FreeSans 100 90 0 0 pix_rst
port 8 ns
<< end >>

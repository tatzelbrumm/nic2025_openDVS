magic
tech sky130A
timestamp 1752335634
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1752335634
transform 1 0 193 0 1 120
box -193 -120 193 120
<< end >>

magic
tech sky130A
timestamp 1752533151
<< isosubstrate >>
rect 0 0 1200 1200
<< metal1 >>
rect 0 944 1200 960
rect 0 976 1200 992
rect 0 1008 1200 1056
rect 0 1072 1200 1096
rect 0 1112 1200 1160
rect 0 1176 1200 1200
<< metal2 >>
rect 1032 0 1056 1200
rect 1072 0 1096 1200
rect 1112 0 1160 1200
rect 1176 0 1200 1200
<< labels >>
flabel metal1 0 1008 1200 1056 0 FreeSans 100 0 0 0 GND
port 0 ew
flabel metal1 0 1112 1200 1160 0 FreeSans 100 0 0 0 VDD
port 1 ew
flabel metal1 0 976 1200 992 0 FreeSans 100 0 0 0 vph_bias
port 2 ew
flabel metal1 0 944 1200 960 0 FreeSans 100 0 0 0 sf_bias
port 3 ew
flabel metal1 0 1072 1200 1096 0 FreeSans 100 0 0 0 vref
port 4 ew
flabel metal1 0 1176 1200 1200 0 FreeSans 100 0 0 0 row_sel
port 5 ew
flabel metal2 1072 0 1096 1200 0 FreeSans 100 90 0 0 sense
port 6 ns
flabel metal2 1032 0 1056 1200 0 FreeSans 100 90 0 0 feedback
port 7 ns
flabel metal2 1176 0 1200 1200 0 FreeSans 100 90 0 0 pix_rst
port 8 ns
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1752622656
<< nmos >>
rect -103 -50 -73 50
rect -15 -50 15 50
rect 73 -50 103 50
<< ndiff >>
rect -161 38 -103 50
rect -161 -38 -149 38
rect -115 -38 -103 38
rect -161 -50 -103 -38
rect -73 38 -15 50
rect -73 -38 -61 38
rect -27 -38 -15 38
rect -73 -50 -15 -38
rect 15 38 73 50
rect 15 -38 27 38
rect 61 -38 73 38
rect 15 -50 73 -38
<< ndiffc >>
rect -149 -38 -115 38
rect -61 -38 -27 38
rect 27 -38 61 38
rect 115 -38 149 38
<< poly >>
rect -103 50 -73 76
rect -15 50 15 76
rect 73 50 103 76
rect -103 -76 -73 -50
rect -15 -76 15 -50
rect 73 -76 103 -50
<< ndiffres >>
rect 103 38 161 50
rect 103 -38 115 38
rect 149 -38 161 38
rect 103 -50 161 -38
<< locali >>
rect -149 38 -115 54
rect -149 -54 -115 -38
rect -61 38 -27 54
rect -61 -54 -27 -38
rect 27 38 61 54
rect 27 -54 61 -38
rect 115 38 149 54
rect 115 -54 149 -38
<< viali >>
rect -149 -38 -115 38
rect -61 -38 -27 38
rect 27 -38 61 38
rect 115 -38 149 38
<< metal1 >>
rect -155 38 -109 50
rect -155 -38 -149 38
rect -115 -38 -109 38
rect -155 -50 -109 -38
rect -67 38 -21 50
rect -67 -38 -61 38
rect -27 -38 -21 38
rect -67 -50 -21 -38
rect 21 38 67 50
rect 21 -38 27 38
rect 61 -38 67 38
rect 21 -50 67 -38
rect 109 38 155 50
rect 109 -38 115 38
rect 149 -38 155 38
rect 109 -50 155 -38
<< end >>

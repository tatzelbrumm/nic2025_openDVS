magic
tech sky130A
timestamp 1752779898
<< isosubstrate >>
rect 0 0 1200 1200
use mimcaps  mimcaps_0
timestamp 1752779898
transform 1 0 187 0 1 448
box 0 0 986 724
use pixeltransistors  pixeltransistors_0
timestamp 1752779898
transform 1 0 760 0 1 580
box 72 -178 377 345
use wires  wires_0
timestamp 1752533151
transform 1 0 0 0 1 0
box 0 0 1200 1200
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1752332266
<< dnwell >>
rect -320 4854 5200 5454
rect -320 534 280 4854
rect 4600 534 5200 4854
rect -320 -66 5200 534
<< photodiode >>
rect 1340 3194 1940 3794
rect 2940 3194 3540 3794
rect 1340 1594 1940 2194
rect 2940 1594 3540 2194
<< nwell >>
rect -400 5248 5280 5534
rect -400 140 -114 5248
rect 1556 3410 1724 3578
rect 3156 3410 3324 3578
rect 1556 1810 1724 1978
rect 3156 1810 3324 1978
rect 4994 140 5280 5248
rect -400 -146 5280 140
<< pwell >>
rect -507 5535 5387 5641
rect -507 -147 -401 5535
rect 5281 -147 5387 5535
rect -507 -253 5387 -147
<< psubdiff >>
rect -471 5571 -375 5605
rect 5255 5571 5351 5605
rect -471 5509 -437 5571
rect 5317 5509 5351 5571
rect -471 -183 -437 -121
rect 5317 -183 5351 -121
rect -471 -217 -375 -183
rect 5255 -217 5351 -183
<< nsubdiff >>
rect -274 5374 -178 5408
rect 5058 5374 5154 5408
rect -274 5312 -240 5374
rect 5120 5312 5154 5374
rect 1599 3511 1681 3535
rect 1599 3477 1623 3511
rect 1657 3477 1681 3511
rect 1599 3453 1681 3477
rect 3199 3511 3281 3535
rect 3199 3477 3223 3511
rect 3257 3477 3281 3511
rect 3199 3453 3281 3477
rect 1599 1911 1681 1935
rect 1599 1877 1623 1911
rect 1657 1877 1681 1911
rect 1599 1853 1681 1877
rect 3199 1911 3281 1935
rect 3199 1877 3223 1911
rect 3257 1877 3281 1911
rect 3199 1853 3281 1877
rect -274 14 -240 76
rect 5120 14 5154 76
rect -274 -20 -178 14
rect 5058 -20 5154 14
<< psubdiffcont >>
rect -375 5571 5255 5605
rect -471 -121 -437 5509
rect 5317 -121 5351 5509
rect -375 -217 5255 -183
<< nsubdiffcont >>
rect -178 5374 5058 5408
rect -274 76 -240 5312
rect 1623 3477 1657 3511
rect 3223 3477 3257 3511
rect 1623 1877 1657 1911
rect 3223 1877 3257 1911
rect 5120 76 5154 5312
rect -178 -20 5058 14
<< locali >>
rect -471 5571 -375 5605
rect 5255 5571 5351 5605
rect -471 5509 -437 5571
rect 5317 5509 5351 5571
rect -274 5374 -178 5408
rect 5058 5374 5154 5408
rect -274 5312 -240 5374
rect 5120 5312 5154 5374
rect 1607 3477 1623 3511
rect 1657 3477 1673 3511
rect 3207 3477 3223 3511
rect 3257 3477 3273 3511
rect 1607 1877 1623 1911
rect 1657 1877 1673 1911
rect 3207 1877 3223 1911
rect 3257 1877 3273 1911
rect -274 14 -240 76
rect 5120 14 5154 76
rect -274 -20 -178 14
rect 5058 -20 5154 14
rect -471 -183 -437 -121
rect 5317 -183 5351 -121
rect -471 -217 -375 -183
rect 5255 -217 5351 -183
<< end >>

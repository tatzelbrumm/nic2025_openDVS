* SPICE3 file created from flatpixels.ext - technology: sky130A

.option scale=5m

D0 a_n471_n217# dw_1340_1594# sky130_fd_pr__model__parasitic__diode_ps2dn area=360000
D1 a_n471_n217# dw_1340_3194# sky130_fd_pr__model__parasitic__diode_ps2dn area=360000
D2 a_n471_n217# dw_2940_1594# sky130_fd_pr__model__parasitic__diode_ps2dn area=360000
D3 a_n471_n217# dw_2940_3194# sky130_fd_pr__model__parasitic__diode_ps2dn area=360000
C0 w_n114_140# dw_n320_n66# 22.2878f
C1 dw_n320_n66# a_n471_n217# 49.4872f

magic
tech sky130A
timestamp 1752857569
<< photodiode >>
rect 0 702 538 790
rect 0 506 630 702
rect 0 364 780 506
rect 0 0 1055 364
<< nwell >>
rect 30 672 508 760
rect 30 476 600 672
rect 30 334 750 476
rect 30 30 1024 334
<< pdiff >>
rect 92 610 445 698
rect 92 414 537 610
rect 92 272 688 414
rect 92 264 957 272
rect 92 100 931 264
rect 948 100 957 264
rect 92 92 957 100
<< pdiffc >>
rect 931 100 948 264
<< psubdiff >>
rect 0 790 17 791
rect 0 773 34 790
rect 504 773 538 790
rect 0 757 17 773
rect 521 756 538 773
rect 521 702 538 719
rect 521 685 555 702
rect 596 685 630 702
rect 613 668 630 685
rect 613 506 630 523
rect 613 489 647 506
rect 746 489 780 506
rect 763 364 780 489
rect 763 347 1054 364
rect 1037 330 1054 347
rect 0 17 17 34
rect 1037 17 1054 34
rect 0 0 34 17
rect 1021 0 1054 17
<< nsubdiff >>
rect 48 725 82 742
rect 456 725 490 742
rect 48 708 65 725
rect 473 708 490 725
rect 473 654 490 671
rect 473 637 507 654
rect 548 637 582 654
rect 565 458 582 475
rect 565 441 599 458
rect 698 441 732 458
rect 715 424 732 441
rect 715 299 732 333
rect 972 299 1006 316
rect 989 282 1006 299
rect 48 65 65 82
rect 989 65 1006 82
rect 48 48 82 65
rect 972 48 1006 65
<< psubdiffcont >>
rect 34 773 504 790
rect 0 34 17 757
rect 521 719 538 756
rect 555 685 596 702
rect 613 523 630 668
rect 647 489 746 506
rect 1037 34 1054 330
rect 34 0 1021 17
<< nsubdiffcont >>
rect 82 725 456 742
rect 48 82 65 708
rect 473 671 490 708
rect 507 637 548 654
rect 565 475 582 637
rect 599 441 698 458
rect 715 333 732 424
rect 732 299 972 316
rect 989 82 1006 282
rect 82 48 972 65
<< locali >>
rect 0 790 17 791
rect 0 773 34 790
rect 504 773 538 790
rect 0 757 17 773
rect 521 756 538 773
rect 48 725 82 742
rect 456 725 490 742
rect 48 708 65 725
rect 473 708 490 725
rect 521 702 538 719
rect 521 685 555 702
rect 596 685 630 702
rect 473 654 490 671
rect 613 668 630 685
rect 473 637 507 654
rect 548 637 582 654
rect 613 506 630 523
rect 613 489 647 506
rect 746 489 780 506
rect 565 458 582 475
rect 565 441 599 458
rect 698 441 732 458
rect 715 424 732 441
rect 763 364 780 489
rect 763 347 1054 364
rect 715 299 732 333
rect 1037 330 1054 347
rect 972 299 1006 316
rect 989 282 1006 299
rect 931 264 948 272
rect 931 92 948 100
rect 48 65 65 82
rect 989 65 1006 82
rect 48 48 82 65
rect 972 48 1006 65
rect 0 17 17 34
rect 1037 17 1054 34
rect 0 0 34 17
rect 1021 0 1054 17
<< labels >>
flabel locali s 931 100 948 264 0 FreeSans 320 90 0 0 anode
port 2 nsew
flabel locali s 82 48 972 65 0 FreeSans 320 0 0 0 cathode
port 1 nsew
flabel locali s 34 0 1021 17 0 FreeSans 320 0 0 0 guard
port 0 nsew
<< end >>

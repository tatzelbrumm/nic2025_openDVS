magic
tech sky130A
magscale 1 2
timestamp 1752626262
<< nmos >>
rect -15 27 15 227
rect -15 -227 15 -27
<< ndiff >>
rect -73 215 -15 227
rect -73 39 -61 215
rect -27 39 -15 215
rect -73 27 -15 39
rect 15 215 73 227
rect 15 39 27 215
rect 61 39 73 215
rect 15 27 73 39
rect -73 -39 -15 -27
rect -73 -215 -61 -39
rect -27 -215 -15 -39
rect -73 -227 -15 -215
rect 15 -39 73 -27
rect 15 -215 27 -39
rect 61 -215 73 -39
rect 15 -227 73 -215
<< ndiffc >>
rect -61 39 -27 215
rect 27 39 61 215
rect -61 -215 -27 -39
rect 27 -215 61 -39
<< poly >>
rect -15 227 15 253
rect -15 -27 15 27
rect -15 -253 15 -227
<< locali >>
rect -61 215 -27 231
rect -61 23 -27 39
rect 27 215 61 231
rect 27 23 61 39
rect -61 -39 -27 -23
rect -61 -231 -27 -215
rect 27 -39 61 -23
rect 27 -231 61 -215
<< viali >>
rect -61 39 -27 215
rect 27 39 61 215
rect -61 -215 -27 -39
rect 27 -215 61 -39
<< metal1 >>
rect -67 215 -21 227
rect -67 39 -61 215
rect -27 39 -21 215
rect -67 27 -21 39
rect 21 215 67 227
rect 21 39 27 215
rect 61 39 67 215
rect 21 27 67 39
rect -67 -39 -21 -27
rect -67 -215 -61 -39
rect -27 -215 -21 -39
rect -67 -227 -21 -215
rect 21 -39 67 -27
rect 21 -215 27 -39
rect 61 -215 67 -39
rect 21 -227 67 -215
<< end >>

magic
tech sky130A
timestamp 1752792418
<< isosubstrate >>
rect 0 0 1200 1200
<< poly >>
rect 1075 985 1108 993
rect 1075 968 1083 985
rect 1101 968 1108 985
rect 1075 960 1108 968
rect 1093 874 1108 960
rect 851 684 884 692
rect 851 667 859 684
rect 876 667 884 684
rect 851 659 884 667
rect 931 684 964 692
rect 931 667 939 684
rect 956 667 964 684
rect 931 659 964 667
rect 861 615 876 659
rect 949 615 964 659
<< polycont >>
rect 1083 968 1101 985
rect 859 667 876 684
rect 939 667 956 684
<< locali >>
rect 1083 1197 1101 1200
rect 1083 985 1101 1177
rect 859 981 876 984
rect 859 684 876 961
rect 1083 960 1101 968
rect 928 939 946 942
rect 928 684 946 919
rect 1114 867 1195 876
rect 1114 781 1177 867
rect 1114 772 1195 781
rect 928 667 939 684
rect 956 667 964 684
rect 859 659 876 667
<< viali >>
rect 1083 1177 1101 1197
rect 859 961 876 981
rect 928 919 946 939
rect 1177 781 1195 867
<< metal1 >>
rect 967 868 1050 874
rect 967 780 1024 868
rect 967 774 1050 780
rect 1174 867 1200 873
rect 1174 775 1200 781
rect 1066 741 1134 747
rect 874 685 907 694
rect 874 659 877 685
rect 904 659 907 685
rect 874 649 907 659
rect 1092 653 1134 741
rect 879 565 902 649
rect 1066 647 1134 653
rect 1023 609 1158 615
rect 1023 421 1108 609
rect 1023 415 1158 421
<< via1 >>
rect 877 1003 904 1047
rect 1024 780 1050 868
rect 1174 781 1177 867
rect 1177 781 1195 867
rect 1195 781 1200 867
rect 877 659 904 685
rect 1066 653 1092 741
rect 1108 421 1158 609
<< metal2 >>
rect 874 1047 907 1050
rect 874 1003 877 1047
rect 904 1003 907 1047
rect 874 685 907 1003
rect 874 659 877 685
rect 904 659 907 685
rect 874 656 907 659
use mimcaps  mimcaps_0
timestamp 1752792418
transform 1 0 187 0 1 448
box 0 0 986 724
use pixeltransistors  pixeltransistors_0
timestamp 1752791877
transform 1 0 760 0 1 580
box 72 -178 377 345
use wires  wires_0
timestamp 1752781518
transform 1 0 0 0 1 0
box 0 0 1200 1200
<< end >>

magic
tech sky130A
timestamp 1752838096
<< nmos >>
rect 233 194 248 294
rect 333 194 348 294
rect 333 67 348 167
rect 101 -15 116 35
rect 145 -15 160 35
rect 189 -15 204 35
rect 289 -165 304 35
<< ndiff >>
rect 204 288 233 294
rect 204 200 210 288
rect 227 200 233 288
rect 204 194 233 200
rect 248 288 277 294
rect 248 200 254 288
rect 271 200 277 288
rect 248 194 277 200
rect 304 288 333 294
rect 304 200 310 288
rect 327 200 333 288
rect 304 194 333 200
rect 348 288 377 294
rect 348 200 354 288
rect 371 200 377 288
rect 348 194 377 200
rect 304 161 333 167
rect 304 73 310 161
rect 327 73 333 161
rect 304 67 333 73
rect 348 161 377 167
rect 348 73 354 161
rect 371 73 377 161
rect 348 67 377 73
rect 72 29 101 35
rect 72 -9 78 29
rect 95 -9 101 29
rect 72 -15 101 -9
rect 116 29 145 35
rect 116 -9 122 29
rect 139 -9 145 29
rect 116 -15 145 -9
rect 160 29 189 35
rect 160 -9 166 29
rect 183 -9 189 29
rect 160 -15 189 -9
rect 260 29 289 35
rect 260 -159 266 29
rect 283 -159 289 29
rect 260 -165 289 -159
rect 304 29 333 35
rect 304 -159 310 29
rect 327 -159 333 29
rect 304 -165 333 -159
<< ndiffc >>
rect 210 200 227 288
rect 254 200 271 288
rect 310 200 327 288
rect 354 200 371 288
rect 310 73 327 161
rect 354 73 371 161
rect 78 -9 95 29
rect 122 -9 139 29
rect 166 -9 183 29
rect 210 -9 227 29
rect 266 -159 283 29
rect 310 -159 327 29
<< psubdiff >>
rect 133 404 421 421
rect 133 146 150 404
rect 28 129 150 146
rect 28 -88 45 129
rect 404 39 421 404
rect 28 -105 168 -88
rect 151 -216 168 -105
rect 360 22 421 39
rect 360 -216 377 22
rect 151 -233 377 -216
<< poly >>
rect 233 337 279 345
rect 233 320 254 337
rect 271 320 279 337
rect 233 312 279 320
rect 233 294 248 312
rect 333 294 348 307
rect 233 181 248 194
rect 333 167 348 194
rect 246 79 279 87
rect 246 62 254 79
rect 271 62 279 79
rect 246 58 279 62
rect 101 35 116 48
rect 145 35 160 48
rect 189 35 204 48
rect 246 43 304 58
rect 333 54 348 67
rect 289 35 304 43
rect 101 -28 116 -15
rect 145 -35 160 -15
rect 189 -28 204 -15
rect 136 -43 169 -35
rect 136 -60 144 -43
rect 161 -60 169 -43
rect 136 -68 169 -60
rect 289 -178 304 -165
<< polycont >>
rect 254 320 271 337
rect 254 62 271 79
rect 144 -60 161 -43
<< ndiffres >>
rect 204 29 233 35
rect 204 -9 210 29
rect 227 -9 233 29
rect 204 -15 233 -9
<< locali >>
rect 133 404 304 421
rect 360 404 421 421
rect 28 129 80 146
rect 133 129 150 404
rect 246 320 254 337
rect 271 320 327 337
rect 210 288 227 296
rect 210 192 227 200
rect 254 288 271 296
rect 28 -88 45 129
rect 254 79 271 200
rect 310 288 327 320
rect 404 314 421 404
rect 310 192 327 200
rect 354 288 371 296
rect 354 192 371 200
rect 254 54 271 62
rect 310 161 327 169
rect 78 29 95 37
rect 78 -43 95 -9
rect 122 29 139 37
rect 122 -17 139 -9
rect 166 29 183 37
rect 166 -17 183 -9
rect 210 29 283 37
rect 227 -9 266 29
rect 210 -17 266 -9
rect 78 -60 144 -43
rect 161 -60 169 -43
rect 28 -105 168 -88
rect 151 -216 168 -105
rect 266 -167 283 -159
rect 310 29 327 73
rect 354 161 371 169
rect 354 65 371 73
rect 404 39 421 173
rect 310 -167 327 -159
rect 360 22 421 39
rect 360 -216 377 22
rect 151 -233 377 -216
<< viali >>
rect 210 200 227 288
rect 78 -9 95 29
rect 122 -9 139 29
rect 166 -9 183 29
rect 210 -9 227 29
rect 266 -159 283 29
rect 354 73 371 161
<< metal1 >>
rect 207 288 230 294
rect 207 200 210 288
rect 227 200 230 288
rect 207 194 230 200
rect 351 161 374 167
rect 351 73 354 161
rect 371 73 374 161
rect 351 67 374 73
rect 75 29 98 35
rect 75 -9 78 29
rect 95 -9 98 29
rect 75 -15 98 -9
rect 119 29 142 35
rect 119 -9 122 29
rect 139 -9 142 29
rect 119 -15 142 -9
rect 163 29 186 35
rect 163 -9 166 29
rect 183 -9 186 29
rect 163 -15 186 -9
rect 207 29 286 35
rect 207 -9 210 29
rect 227 -9 266 29
rect 207 -15 266 -9
rect 263 -159 266 -15
rect 283 -159 286 29
rect 263 -165 286 -159
<< end >>

magic
tech sky130A
timestamp 1752840811
<< error_s >>
rect 903 347 1037 360
<< poly >>
rect 1075 959 1108 967
rect 1075 942 1083 959
rect 1101 942 1108 959
rect 1075 934 1108 942
rect 1093 874 1108 934
rect 851 684 884 692
rect 851 667 859 684
rect 876 667 884 684
rect 851 659 884 667
rect 931 684 964 692
rect 931 667 939 684
rect 956 667 964 684
rect 931 659 964 667
rect 861 615 876 659
rect 949 615 964 659
rect 944 407 977 415
rect 944 390 952 407
rect 969 399 977 407
rect 1049 399 1064 415
rect 969 390 1064 399
rect 944 382 1064 390
<< polycont >>
rect 1083 942 1101 959
rect 859 667 876 684
rect 939 667 956 684
rect 952 390 969 407
<< locali >>
rect 1083 1197 1101 1200
rect 859 981 876 984
rect 859 684 876 961
rect 1083 959 1101 1177
rect 928 939 946 942
rect 1083 934 1101 942
rect 928 684 946 919
rect 1114 867 1195 876
rect 1114 781 1177 867
rect 1114 772 1195 781
rect 928 667 939 684
rect 956 667 964 684
rect 859 659 876 667
rect 944 407 977 415
rect 944 390 952 407
rect 969 390 977 407
rect 944 382 977 390
<< viali >>
rect 1083 1177 1101 1197
rect 859 961 876 981
rect 928 919 946 939
rect 1177 781 1195 867
rect 1120 421 1137 602
rect 952 390 969 407
<< metal1 >>
rect 967 868 1050 874
rect 967 780 1024 868
rect 967 774 1050 780
rect 1174 867 1200 873
rect 1174 775 1200 781
rect 1066 741 1134 747
rect 515 710 946 733
rect 515 708 554 710
rect 515 681 521 708
rect 548 681 554 708
rect 515 675 554 681
rect 874 685 907 694
rect 874 659 877 685
rect 904 659 907 685
rect 874 649 907 659
rect 879 565 902 649
rect 923 565 946 710
rect 1092 653 1134 741
rect 1066 647 1134 653
rect 1023 609 1158 615
rect 1023 421 1108 609
rect 1023 415 1158 421
rect 944 412 977 415
rect 944 385 947 412
rect 974 385 977 412
rect 944 382 977 385
<< via1 >>
rect 761 1066 792 1092
rect 877 1003 904 1047
rect 1024 780 1050 868
rect 1174 781 1177 867
rect 1177 781 1195 867
rect 1195 781 1200 867
rect 521 681 548 708
rect 877 659 904 685
rect 1066 653 1092 741
rect 1108 602 1158 609
rect 1108 421 1120 602
rect 1120 421 1137 602
rect 1137 421 1158 602
rect 947 407 974 412
rect 947 390 952 407
rect 952 390 969 407
rect 969 390 974 407
rect 947 385 974 390
<< metal2 >>
rect 759 1092 794 1095
rect 759 1066 761 1092
rect 792 1066 794 1092
rect 515 709 554 714
rect 515 680 520 709
rect 549 680 554 709
rect 515 675 554 680
rect 759 418 794 1066
rect 874 1047 907 1050
rect 874 1003 877 1047
rect 904 1003 907 1047
rect 874 685 907 1003
rect 874 659 877 685
rect 904 659 907 685
rect 874 656 907 659
rect 757 413 796 418
rect 757 384 762 413
rect 791 384 796 413
rect 757 379 796 384
rect 936 413 984 424
rect 936 384 946 413
rect 975 384 984 413
rect 936 376 984 384
<< via2 >>
rect 520 708 549 709
rect 520 681 521 708
rect 521 681 548 708
rect 548 681 549 708
rect 520 680 549 681
rect 762 384 791 413
rect 946 412 975 413
rect 946 385 947 412
rect 947 385 974 412
rect 974 385 975 412
rect 946 384 975 385
<< metal3 >>
rect 508 712 560 720
rect 508 678 517 712
rect 552 678 560 712
rect 508 672 560 678
rect 750 416 802 424
rect 750 382 759 416
rect 794 382 802 416
rect 750 376 802 382
rect 934 416 986 424
rect 934 382 943 416
rect 978 382 986 416
rect 934 376 986 382
<< via3 >>
rect 517 709 552 712
rect 517 680 520 709
rect 520 680 549 709
rect 549 680 552 709
rect 517 678 552 680
rect 759 413 794 416
rect 759 384 762 413
rect 762 384 791 413
rect 791 384 794 413
rect 759 382 794 384
rect 943 413 978 416
rect 943 384 946 413
rect 946 384 975 413
rect 975 384 978 413
rect 943 382 978 384
<< metal4 >>
rect 510 712 558 833
rect 510 678 517 712
rect 552 678 558 712
rect 510 672 558 678
rect 752 416 800 536
rect 752 382 759 416
rect 794 382 800 416
rect 752 376 800 382
rect 936 416 984 482
rect 936 382 943 416
rect 978 382 984 416
rect 936 376 984 382
use mimcaps  mimcaps_0
timestamp 1752840811
transform 1 0 0 0 1 476
box 0 0 986 724
use photodiode  photodiode_0
timestamp 1752840811
transform 1 0 0 0 1 0
box 0 0 1024 760
use pixeltransistors  pixeltransistors_0
timestamp 1752839314
transform 1 0 760 0 1 580
box 28 -233 421 421
use wires  wires_0
timestamp 1752839314
transform 1 0 0 0 1 0
box 0 0 1200 1200
<< end >>
